// WSA1000 is receive-only.
`include "../include/common_config_2rxhb_0tx.vh"

`include "../include/common_config_bottom.vh"
